
module lab62_soc (
	acc_wire_export,
	clk_clk,
	hex_digits_export,
	i2c_wire_sda_in,
	i2c_wire_scl_in,
	i2c_wire_sda_oe,
	i2c_wire_scl_oe,
	key0_wire_export,
	key1_wire_export,
	key_external_connection_export,
	keycode_export,
	leds_export,
	reset_reset_n,
	sdram_clk_clk,
	sdram_wire_addr,
	sdram_wire_ba,
	sdram_wire_cas_n,
	sdram_wire_cke,
	sdram_wire_cs_n,
	sdram_wire_dq,
	sdram_wire_dqm,
	sdram_wire_ras_n,
	sdram_wire_we_n,
	spi0_MISO,
	spi0_MOSI,
	spi0_SCLK,
	spi0_SS_n,
	sw_wire_export,
	usb_gpx_export,
	usb_irq_export,
	usb_rst_export,
	vga_port_red,
	vga_port_green,
	vga_port_blue,
	vga_port_hs,
	vga_port_vs);	

	input		acc_wire_export;
	input		clk_clk;
	output	[15:0]	hex_digits_export;
	input		i2c_wire_sda_in;
	input		i2c_wire_scl_in;
	output		i2c_wire_sda_oe;
	output		i2c_wire_scl_oe;
	input		key0_wire_export;
	input		key1_wire_export;
	input	[1:0]	key_external_connection_export;
	output	[7:0]	keycode_export;
	output	[13:0]	leds_export;
	input		reset_reset_n;
	output		sdram_clk_clk;
	output	[12:0]	sdram_wire_addr;
	output	[1:0]	sdram_wire_ba;
	output		sdram_wire_cas_n;
	output		sdram_wire_cke;
	output		sdram_wire_cs_n;
	inout	[15:0]	sdram_wire_dq;
	output	[1:0]	sdram_wire_dqm;
	output		sdram_wire_ras_n;
	output		sdram_wire_we_n;
	input		spi0_MISO;
	output		spi0_MOSI;
	output		spi0_SCLK;
	output		spi0_SS_n;
	input	[9:0]	sw_wire_export;
	input		usb_gpx_export;
	input		usb_irq_export;
	output		usb_rst_export;
	output	[3:0]	vga_port_red;
	output	[3:0]	vga_port_green;
	output	[3:0]	vga_port_blue;
	output		vga_port_hs;
	output		vga_port_vs;
endmodule
